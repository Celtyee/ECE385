module BEN_Unit(
    input logic Clk, Reset
);