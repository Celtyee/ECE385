module datapath (
    input logic[15:0] Gate_MAR, Gate_PC, Gate_MDR, Gate_ALU,
    input logic[3:0] choose_sig,
    output logic[15:0] data
);
    case(choose_sig)
    
endmodule