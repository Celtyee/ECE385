    Mac OS X            	   2  �     �                                    ATTR     �   �   I                  �   9  com.apple.quarantine    �     com.apple.lastuseddate#PS 9E-0083;5e610a86;Safari;65E5CC80-1505-4E9E-80B9-95A5F4E856FA`N{^    �x�*                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          This resource fork intentionally left blank                                                                                                                                                                                                                            ��