// 1
module Instruction_adder (
    input logic [15:0]
);
    
endmodule

//2
module IR (
    ports
);
    
endmodule

//3
module BR_logic (
    ports
);
    
endmodule

//4
module REG_FILE (
    ports
);
    
endmodule

//5
module PC_Count (
    ports
);
    
endmodule

//6
module ALUK (
    ports
);
    
endmodule

//7
module ALU (
    ports
);
    
endmodule
