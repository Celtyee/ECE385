module REG_FILE (
    input logic Clk, Reset_ah, DR, SR1, LD_REG,
    input logic [15:0] datapath_out,
    input logic [2:0] IR_11_9, IR_8_6,SR2,
    output logic [15:0] SR1_out, SR2_out
);
    
endmodule

