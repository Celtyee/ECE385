    Mac OS X            	   2  �     �                                    ATTR     �   �  E                  �   9  com.apple.quarantine       %com.apple.metadata:kMDItemWhereFroms 0081;5e7861e2;Chrome;117B97BB-A840-4FB1-89D7-F98B681601BFbplist00�_rhttps://c.zju.edu.cn/bbcswebdav/pid-142845-dt-content-rid-3403429_1/courses/UIUC-1001921-h117043-3668/testbench.sv_fhttps://c.zju.edu.cn/webapps/blackboard/content/listContent.jsp?course_id=_5268_1&content_id=_133644_1�                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  This resource fork intentionally left blank                                                                                                                                                                                                                            ��