module IR_ADDER #(W=16)(
    input logic Clk, Reset_ah,
    output logic [W-1:0] adder_output
);
    
endmodule